library IEEE;
use IEEE.STD_Logic_1164.all;
USE ieee.numeric_std.ALL; 

entity print is
	PORT(
		clk_vga					:	in STD_LOGIC;
		column, row				:	in INTEGER;
		vga_R, vga_G,vga_B	:	out STD_LOGIC_VECTOR(3 downto 0);
		pintar					:	in	STD_LOGIC;
		L, R, U, D				:	in STD_LOGIC;
		shoot						:  in STD_LOGIC;
		btnB						:	in std_logic
	);
end;
 
architecture behavioral of print is


--------------------------------------------
--------------- Componentes ----------------
--------------------------------------------

component random is
	Port (
			clk : in STD_LOGIC;
			en : in STD_LOGIC;
			random_number : out STD_LOGIC_VECTOR (8 downto 0)
	);
end component;

component divisorPrint is
	Port (
			clk_vga : in STD_LOGIC;
			clk25   : out STD_LOGIC
	);
end component;
--

--------------------------------------------
---------------- Constantes ----------------
--------------------------------------------

-- Resolucion de la imagen de salida
constant h_video	:	INTEGER := 640;	-- pixeles horizontales
constant v_video	:	INTEGER := 480;	-- pixeles verticales
constant tam		:	INTEGER := 30;		-- Tamaño de la nave 30x30
constant radio_asteroide : INTEGER := 10;
constant distancia : INTEGER := 60;		-- distancia vertical entre cada asteroide
constant tam_disp : INTEGER := 10;	-- Tamaño del disparo

-----------------------------------------------
----------------- Mapas de bits ---------------
-----------------------------------------------
											
type imagen30 is array (0 to 899) of STD_LOGIC_vector(11 downto 0);
constant vector_nave : imagen30 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"000",x"000",x"000",x"000",x"100",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"001",x"001",x"001",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"012",x"123",x"123",x"012",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"112",x"123",x"123",x"012",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"112",x"123",x"123",x"012",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"112",x"123",x"123",x"012",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"112",x"123",x"123",x"112",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"211",x"322",x"322",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"211",x"321",x"321",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"211",x"211",x"221",x"321",x"321",x"221",x"211",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"321",x"321",x"321",x"331",x"331",x"321",x"321",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"321",x"321",x"321",x"331",x"331",x"321",x"321",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"321",x"321",x"321",x"331",x"331",x"321",x"321",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"321",x"321",x"321",x"331",x"331",x"321",x"321",x"311",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"112",x"112",x"012",x"000",x"100",x"321",x"321",x"321",x"331",x"331",x"321",x"321",x"211",x"000",x"000",x"012",x"112",x"012",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"001",x"123",x"123",x"122",x"000",x"100",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"000",x"001",x"123",x"123",x"123",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"001",x"123",x"123",x"122",x"100",x"100",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"000",x"101",x"123",x"123",x"123",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"001",x"123",x"123",x"222",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"311",x"211",x"211",x"123",x"123",x"122",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"001",x"123",x"123",x"223",x"211",x"311",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"223",x"123",x"123",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"110",x"211",x"211",x"222",x"223",x"222",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"222",x"223",x"222",x"211",x"211",x"100",x"000",x"000",x"000",
	x"000",x"000",x"000",x"211",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"211",x"000",x"000",x"000",
	x"000",x"100",x"100",x"211",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"211",x"100",x"100",x"000",
	x"100",x"311",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"311",x"311",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"000",
	x"110",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"000",
	x"110",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"311",x"100",
	x"100",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"311",x"100",
	x"100",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"321",x"321",x"321",x"321",x"321",x"311",x"000",
	x"100",x"211",x"211",x"211",x"211",x"211",x"211",x"211",x"211",x"110",x"211",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"311",x"110",x"110",x"211",x"211",x"211",x"211",x"211",x"211",x"211",x"211",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"321",x"321",x"321",x"211",x"211",x"321",x"321",x"311",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"211",x"321",x"211",x"211",x"211",x"311",x"321",x"211",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
--

type imagen100 is array (0 to 9999) of STD_LOGIC_vector(11 downto 0);
constant vector_over : imagen100 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"EEE",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"EEE",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"EEE",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",x"000",x"000",x"000",x"EEE",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"EEE",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
	
--

type number24 is array (0 to 575) of std_logic_vector(11 downto 0);
constant numero0 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);

constant numero1 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero2 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero3 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero4 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero5 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero6 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero7 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero8 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
constant numero9 : number24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
--

type corazon24 is array (0 to 575) of STD_LOGIC_vector(11 downto 0); 
constant cora : corazon24 := 
(
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"FFF",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",
	x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"FFF",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",
	x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",
	x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",
	x"000",x"000",x"000",x"FFF",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"F00",x"F00",x"F00",x"F00",x"F00",x"F00",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"F00",x"F00",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
	x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"FFF",x"FFF",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"
);
--


-----------------------------------------------
------------------ Señales --------------------
-----------------------------------------------

--- Desplazamiento en X y Y para mover la nave
signal despX	: INTEGER range -1 to 640:=305; -- Valores iniciales para posicionar la nave justo en el centro de la
signal despY	: INTEGER range -1 to 480:= v_video-tam-1; -- parte inferior de la pantalla cuando se inicia el juego

-- Definimos las señales que nos inidicaran el desplazamiento en Y de los asteroides
-- Esta desplazamiento está dado por la señal de reloj de 25 Hz
signal desp_asteroide0 : integer range -1 to 480 := 0;
signal desp_asteroide1 : integer range -1 to 480 := 0;
signal desp_asteroide2 : integer range -1 to 480 := 0;
signal desp_asteroide3 : integer range -1 to 480 := 0;
signal desp_asteroide4 : integer range -1 to 480 := 0;
signal desp_asteroide5 : integer range -1 to 480 := 0;
signal desp_asteroide6 : integer range -1 to 480 := 0;
signal desp_asteroide7 : integer range -1 to 480 := 0;

-- Posicion en X de los asteroides, que será aleaotoria
signal posX_asteroide0 : integer range 0 to 640 := 0;
signal posX_asteroide1 : integer range 0 to 640 := 0;
signal posX_asteroide2 : integer range 0 to 640 := 0;
signal posX_asteroide3 : integer range 0 to 640 := 0;
signal posX_asteroide4 : integer range 0 to 640 := 0;
signal posX_asteroide5 : integer range 0 to 640 := 0;
signal posX_asteroide6 : integer range 0 to 640 := 0;
signal posX_asteroide7 : integer range 0 to 640 := 0;
-- posX_asteroide y desp_asteroide, serán las coordenadas del centro de cada asteroide

-- Desplazamiento en Y del disparo
signal desp_disparo	  : INTEGER range -1 to 480:=470;
-- Posicion en X del disparo
signal posx_disparo    : integer range 0 to 640 := 0;
-- disparo activo
signal recarga         : std_logic := '1';

--- Banderas que nos indican si los contadores en X e Y entran en el rango válido
-- de cada uno de los elementos. Ya sea la nave o el asteroide
signal nave_vali	: std_logic := '0';
signal ast_vali0	: std_logic := '0';
signal ast_vali1	: std_logic := '0';
signal ast_vali2	: std_logic := '0';
signal ast_vali3	: std_logic := '0';
signal ast_vali4	: std_logic := '0';
signal ast_vali5	: std_logic := '0';
signal ast_vali6	: std_logic := '0';
signal ast_vali7	: std_logic := '0';
signal disparo_vali: std_logic := '0';


--- Banderas de explosion
signal explota_asteroide0, explota_asteroide1, explota_asteroide2, explota_asteroide3 : std_logic := '0'; 
signal explota_asteroide4, explota_asteroide5, explota_asteroide6, explota_asteroide7 : std_logic := '0';
signal explota_disparo : std_logic := '0';
signal explota_nave : std_logic := '0';

-- Este ultimo es para hacer un OR con todas las anteriores ya que sólo basta con que
-- una de las banderas de los asteroides se active para mandar la señal del color al vga
signal asteroide_valido	: std_logic := '0';
signal vel_asteroide : integer range 0 to 7 := 0;

--- Señal de reloj a 25H para el movimiento de la nave y asteroides
signal clk25	: STD_LOGIC := '0';

-- Señal que se le envía al VGA
signal vga_color : STD_LOGIC_VECTOR(11 downto 0):= x"000";

-- Color de cada pixel de que define a los objetos
signal color_nave : STD_LOGIC_VECTOR(11 downto 0) := x"000";
signal color_over : STD_LOGIC_VECTOR(11 downto 0) := x"000";
signal color_numero1 : std_logic_vector(11 downto 0) := x"000";
signal color_numero2 : std_logic_vector(11 downto 0) := x"000";
signal color_numero3 : std_logic_vector(11 downto 0) := x"000";
signal color_cora1	: std_logic_vector(11 downto 0) := x"000";
signal color_cora2	: std_logic_vector(11 downto 0) := x"000";
signal color_cora3	: std_logic_vector(11 downto 0) := x"000";

signal over_vali : std_logic := '0';
-- Banderas para los digitos del contador
signal num1_vali : std_logic := '0';
signal num2_vali : std_logic := '0';
signal num3_vali : std_logic := '0';
-- Banderas para las vidas disponibles
signal cor1_vali : std_logic := '0';
signal cor2_vali : std_logic := '0';
signal cor3_vali : std_logic := '0';

-- Seña de start para inciar el juego
signal start : std_logic := '0';

-- Contador de asteroides destruidos
signal destruidos : integer range 0 to 1000 := 0;

-- Contador de vidas
signal vidas : integer range 0 to 3 := 3;
signal reiniciar : std_logic := '0';

-- Numero Random para la posicion en x de los asteroides
signal numero_random : std_logic_vector (8 downto 0);
shared variable gen_random		: std_logic := '0';  -- Bandera que se activa cuando se quiere generar un numero random
																	-- Es de tipo variable para que cambia su valor al instante y no se espere
																	-- hasta que finalice el proceso, de esta manera se genera el numero random
																	-- de manera inmediata

------------------------------------------------------
------------------- Procesos -------------------------
------------------------------------------------------																	
																
begin
	
	-- Mapeamos nuestra entiendad 
	generar_random : random port map(clk_vga,gen_random,numero_random);

	-- Divisor de frecuencia a 25 Hz 
	divisor_25 : divisorPrint port map(clk_vga, clk25);
	
	-- Proceso para iniciar al juego
	iniciar : process (clk_vga, vidas) is
	begin 
		if rising_edge(clk_vga) then
			if btnB = '1' then
				start <= '1';
			elsif vidas = 0 then
				start <= '0';
			end if;
		end if;
	end process iniciar;
	--
	
	quitar_vida : process (explota_nave)
	begin
		if explota_nave = '1' then
			vidas <= vidas-1;
		end if;
	end process quitar_vida;
	--
	
	-- Este proceso Aumenta o decrementa los contadores en X e Y que definen el rango en el cual se mostrará la nave.
	mover_nave : process (clk25,L,R, U,D) is 
	begin
		if rising_edge(clk25) then
			if start = '1' then
				if L = '1' then
					despX <= despX - 1;
				end if;
				if R = '1' then
					despX <= despX + 1;
				end if;
				
				if U = '1' then
					despY <= despY - 1;
				end if;
				if D = '1' then
					despY <= despY + 1;
				end if;
				
				-- Bordes
				if despX = h_video-tam-111 then
					despX <= h_video-tam-112;
				elsif despX = 0 then
					despX <= 1;
				end if;
				
				if despY = v_video-tam-1 then
					despY <= v_video-tam-2;
				elsif despY = 0 then
					despY <= 1;
				end if;
			else
				despX	<=305;
				despY	<=v_video-tam-1;
			end if;
		end if;
	end process mover_nave;
	--
	
	disparar : process(clk25, shoot, recarga, explota_disparo, desp_disparo) is
		--- Proceso para iniciar el disparo, si recarga es = 0 entonces dispara, ya que no hay un disparo
		--- activo, si es = 1, no pasa nada. Cuando se dispara se cambia el estado a activado y se asigna el 
		--- valor de x donde se genera el disparo
	begin		
		if rising_edge(clk25) then
			if start = '1' then
				if explota_disparo = '1' then
					desp_disparo <= despY;
					recarga <= '1';
					
				else
					-- validacion de disparo
					if recarga = '1' then
						if shoot = '1' then
							posx_disparo <= despx + 15 - tam_disp/2; -- dispara en donde empieza + nave a la mitad
							desp_disparo <= despY;
							recarga <= '0';
						end if;
					else
					--	--- Mueve el cuadrito del disparo
						if desp_disparo > 0 then
							desp_disparo <= desp_disparo-5;
							recarga <= '0';
						else
							desp_disparo <= despY;
							recarga <= '1';
						end if;
					end if;
				end if;
			else
				desp_disparo <= despY;
				recarga <= '1';
			end if;
		end if;
	end process disparar;
	--
	
	-- Este proces detecta la colision de algun asteroide con la nave
	impacto_nave : process (clk25, U) is
	begin
		if rising_edge(clk25) then
			if desp_asteroide0+radio_asteroide > 450 and desp_asteroide0+radio_asteroide < 479 and
				despX > posX_asteroide0-radio_asteroide-30 and despX < posX_asteroide0+radio_asteroide then
				explota_nave  <= '1';
				
			elsif desp_asteroide1+radio_asteroide > 450 and desp_asteroide1+radio_asteroide < 479 and
				despX > posX_asteroide1-radio_asteroide-30 and despX < posX_asteroide1+radio_asteroide then
				explota_nave  <= '1';
			
			elsif desp_asteroide2+radio_asteroide > 450 and desp_asteroide2+radio_asteroide < 479 and
				despX > posX_asteroide2-radio_asteroide-30 and despX < posX_asteroide2+radio_asteroide then
				explota_nave  <= '1';
				
			elsif desp_asteroide2+radio_asteroide > 450 and desp_asteroide2+radio_asteroide < 479 and
				despX > posX_asteroide2-radio_asteroide-30 and despX < posX_asteroide2+radio_asteroide then
				explota_nave  <= '1';
			
			elsif desp_asteroide3+radio_asteroide > 450 and desp_asteroide3+radio_asteroide < 479 and
				despX > posX_asteroide3-radio_asteroide-30 and despX < posX_asteroide3+radio_asteroide then
				explota_nave  <= '1';
			
			elsif desp_asteroide4+radio_asteroide > 450 and desp_asteroide4+radio_asteroide < 479 and
				despX > posX_asteroide4-radio_asteroide-30 and despX < posX_asteroide4+radio_asteroide then
				explota_nave  <= '1';
				
			elsif desp_asteroide5+radio_asteroide > 450 and desp_asteroide5+radio_asteroide < 479 and
				despX > posX_asteroide5-radio_asteroide-30 and despX < posX_asteroide5+radio_asteroide then
				explota_nave  <= '1';
				
			elsif desp_asteroide6+radio_asteroide > 450 and desp_asteroide6+radio_asteroide < 479 and
				despX > posX_asteroide6-radio_asteroide-30 and despX < posX_asteroide6+radio_asteroide then
				explota_nave  <= '1';
				
			elsif desp_asteroide7+radio_asteroide > 450 and desp_asteroide7+radio_asteroide < 479 and
				despX > posX_asteroide7-radio_asteroide-30 and despX < posX_asteroide7+radio_asteroide then
				explota_nave  <= '1';
			
			else
				if start = '1' then
					explota_nave <= '0';
				end if;
			end if;
				
		end if;
		
	end process impacto_nave;
	--
	
	-- Este proceso detecta cuando un disparo choca con algun asteroide.
	impacto_asteroide : process(clk25) is
	begin
		if rising_edge(clk25) then
			if vidas = 0 and btnB = '1' then
				destruidos <= 0;
			end if;
			
			if recarga = '0' then
				if desp_disparo < desp_asteroide0+radio_asteroide
					and posx_disparo > posX_asteroide0-radio_asteroide-10 and posx_disparo < posX_asteroide0+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide0 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide1+radio_asteroide
					and posx_disparo > posX_asteroide1-radio_asteroide-10 and posx_disparo < posX_asteroide1+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide1 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide2+radio_asteroide 
					and posx_disparo > posX_asteroide2-radio_asteroide-10 and posx_disparo < posX_asteroide2+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide2 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide3+radio_asteroide
					and posx_disparo > posX_asteroide3-radio_asteroide-10 and posx_disparo < posX_asteroide3+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide3 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide4+radio_asteroide
					and posx_disparo > posX_asteroide4-radio_asteroide-10 and posx_disparo < posX_asteroide4+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide4 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide5+radio_asteroide
					and posx_disparo > posX_asteroide5-radio_asteroide-10 and posx_disparo < posX_asteroide5+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide5 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide6+radio_asteroide 
					and posx_disparo > posX_asteroide6-radio_asteroide-10 and posx_disparo < posX_asteroide6+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide6 <= '1';
					destruidos <= destruidos + 1;
				
				elsif desp_disparo < desp_asteroide7+radio_asteroide
					and posx_disparo > posX_asteroide7-radio_asteroide-10 and posx_disparo < posX_asteroide7+radio_asteroide then
					explota_disparo <= '1';
					explota_asteroide6 <= '1';
					destruidos <= destruidos + 1;
				
				elsif vidas = 0 then
					explota_disparo <= '1';
				end if;
			
			else 
				explota_disparo <= '0';
				explota_asteroide0 <= '0';
				explota_asteroide1 <= '0';
				explota_asteroide2 <= '0';
				explota_asteroide3 <= '0';
				explota_asteroide4 <= '0';
				explota_asteroide5 <= '0';
				explota_asteroide6 <= '0';
				explota_asteroide7 <= '0';
			end if;
		
		end if;
		
	end process impacto_asteroide;
	--
	
	--Proceso que posiciona aleatoriamente en X el asteroide cuando este llega hasta abajo
	posicionar_asteroide : process (numero_random,desp_asteroide0,desp_asteroide1,desp_asteroide2,desp_asteroide3,desp_asteroide4,desp_asteroide5,desp_asteroide6,desp_asteroide7) is
	begin
		
		-- Este proceso Detecta cuando el contador en Y (desp_asteroide) de cada asteroide ha llegado hasta
		-- abajo (499), si es así entonces activa la señal para generar un numero aleatorio y lo asigna a la posicion
		-- en X (posX_asteroide) del asteroide en cuestión. Así cuando vuelva a aparecer en la parte superior su posicion
		-- en X será aleatoria
		-- Ocupamos elsif y no if independientes porque los asteroides van un tras otro, entonces
		-- no se puede dar el caso en el que dos o más lleguen al fondo al mismo tiempo, ya que los
		-- contadores en Y de cada uno están desplazados lo que indica la constante 'distancia'
		
		if desp_asteroide0 >= 479 then
			gen_random := '1';
			posX_asteroide0 <= to_integer(unsigned(numero_random));

		elsif desp_asteroide1 >= 479 then
			gen_random := '1';
			posX_asteroide1 <= to_integer(unsigned(numero_random));
		
		elsif desp_asteroide2 >= 479 then
			gen_random := '1';
			posX_asteroide2 <= to_integer(unsigned(numero_random));

		elsif desp_asteroide3 >= 479 then
			gen_random := '1';
			posX_asteroide3 <= to_integer(unsigned(numero_random));

		elsif desp_asteroide4 >= 479 then
			gen_random := '1';
			posX_asteroide4 <= to_integer(unsigned(numero_random));

		elsif desp_asteroide5 >= 479 then
			gen_random := '1';
			posX_asteroide5 <= to_integer(unsigned(numero_random));

		elsif desp_asteroide6 >= 479 then
			gen_random := '1';
			posX_asteroide6 <= to_integer(unsigned(numero_random));

		elsif desp_asteroide7 >= 479 then
			gen_random := '1';
			posX_asteroide7 <= to_integer(unsigned(numero_random));
			
		-- Si ninguno de los asteroides ha llegado al fondo entonces
		-- apagamos la bandera de los numero aleatorios 
		else
			gen_random := '0';
		end if;
		
		
	end process posicionar_asteroide;
	--
	
	velocidad_asteroide: process(clk_vga) is
	begin 
		if rising_edge(clk_vga) then
			if destruidos < 50 then
				vel_asteroide <= 0;
			elsif destruidos >= 50 and destruidos < 100 then
				vel_asteroide <= 1;
			elsif destruidos >= 100 and destruidos < 150 then
				vel_asteroide <= 2;
			elsif destruidos >= 150 and destruidos < 200 then
				vel_asteroide <= 3;
			elsif destruidos >= 200 and destruidos < 250 then
				vel_asteroide <= 4;
			elsif destruidos >= 250 and destruidos < 300 then
				vel_asteroide <= 5;
			elsif destruidos >= 300 and destruidos < 350 then
				vel_asteroide <= 6;
			end if;
		end if;
	end process velocidad_asteroide;
	
	
	
	-- Proceso que aumenta el contador en Y de cada asteroide por cada ciclo de reloj
	mover_asteroide : process(clk25,explota_asteroide0,explota_asteroide1,explota_asteroide2,explota_asteroide3,explota_asteroide4,explota_asteroide5,explota_asteroide6,explota_asteroide7) is
		-- varifica que si se ha llegado al fondo el contador se reinicie. Además, asegura que cada contador
		-- no empiece su cuenta hasta que el contador del asteroide anterior haya llegada a la distancia de
		-- separación que se le indico en la constante 'distancia'
	begin
		
		if rising_edge(clk25) then	
			if start = '1' then
				-- mueve asteroides y aumenta su vellcidad cada 50 puntos
				if desp_asteroide0 >= 479 then
					desp_asteroide0 <= 0;
				elsif explota_asteroide0 = '1' then
					desp_asteroide0 <= 479;
				else
					desp_asteroide0 <= desp_asteroide0+1+vel_asteroide;
				end if;

				if desp_asteroide1 >= 479 or (desp_asteroide0<distancia and desp_asteroide1=0)then
					desp_asteroide1 <= 0;
				elsif explota_asteroide1 = '1' then
					desp_asteroide1 <= 479;
				else
					desp_asteroide1 <= desp_asteroide1+1+vel_asteroide;
				end if;
				
				if desp_asteroide2 >= 479 or (desp_asteroide1<distancia and desp_asteroide2=0) then
					desp_asteroide2 <= 0;
				elsif explota_asteroide2 = '1' then
					desp_asteroide2 <= 479;
				else
					desp_asteroide2 <= desp_asteroide2+1+vel_asteroide;
				end if;

				if desp_asteroide3 >= 479 or (desp_asteroide2<distancia and desp_asteroide3=0) then
					desp_asteroide3 <= 0;
				elsif explota_asteroide3 = '1' then
					desp_asteroide3 <= 479;
				else
					desp_asteroide3 <= desp_asteroide3+1+vel_asteroide;
				end if;

				if desp_asteroide4 >= 479 or (desp_asteroide3<distancia and desp_asteroide4=0) then
					desp_asteroide4 <= 0;
				elsif explota_asteroide4 = '1' then
					desp_asteroide4 <= 479;
				else
					desp_asteroide4 <= desp_asteroide4+1+vel_asteroide;
				end if;

				if desp_asteroide5 >= 479 or (desp_asteroide4<distancia and desp_asteroide5=0) then
					desp_asteroide5 <= 0;
				elsif explota_asteroide5 = '1' then
					desp_asteroide5 <= 479;
				else
					desp_asteroide5 <= desp_asteroide5+1+vel_asteroide;
				end if;

				if desp_asteroide6 >= 479 or (desp_asteroide5<distancia and desp_asteroide6=0) then
					desp_asteroide6 <= 0;
				elsif explota_asteroide6 = '1' then
					desp_asteroide6 <= 479;
				else
					desp_asteroide6 <= desp_asteroide6+1+vel_asteroide;
				end if;

				if desp_asteroide7 >= 479 or (desp_asteroide6<distancia and desp_asteroide7=0) then
					desp_asteroide7 <= 0;
				elsif explota_asteroide7 = '1' then
					desp_asteroide7 <= 479;
				else
					desp_asteroide7 <= desp_asteroide7+1+vel_asteroide;
				end if;
			else
				desp_asteroide0 <= 0;
				desp_asteroide1 <= 0;
				desp_asteroide2 <= 0;
				desp_asteroide3 <= 0;
				desp_asteroide4 <= 0;
				desp_asteroide5 <= 0;
				desp_asteroide6 <= 0;
				desp_asteroide7 <= 0;
				
			end if;
		end if;
	end process mover_asteroide;
	--
	
	-- Contador que nos va idicando en que posicion del arreglo de la nave colocarnos
	contador_nave : process (clk_vga, nave_vali) is
		variable contador : integer range -1 to 900 := -1;
	begin
		if rising_edge(clk_vga) then
			if nave_vali = '1' then
				contador := contador+1;
				if contador = 899 then
					contador := -1;
				end if;
			end if;
		end if;
		color_nave <= vector_nave(contador);
	end process contador_nave;
	--
	
	contador_over : process (clk_vga, over_vali) is
		variable contador : integer range -1 to 10000 := -1;
	begin
		if rising_edge(clk_vga) then
			if over_vali = '1' then
				contador := contador+1;
				if contador = 9999 then
					contador := -1;
				end if;
			end if;
		end if;
		color_over <= vector_over(contador);
	end process contador_over;
	--
	
	contador_numero1 : process (clk_vga, num1_vali) is
		variable contador : integer range -1 to 576 := -1;
	begin	
		if rising_edge(clk_vga) then
			if num1_vali = '1' then
				contador := contador+1;
				if contador = 575 then
					contador := -1;
				end if;
			end if;
		end if;
		
		if destruidos/100 = 0 then
			color_numero1 <= numero0(contador);
		elsif destruidos/100 = 1 then
			color_numero1 <= numero1(contador);
		elsif destruidos/100 = 2 then
			color_numero1 <= numero2(contador);
		elsif destruidos/100 = 3 then
			color_numero1 <= numero3(contador);
		elsif destruidos/100 = 4 then
			color_numero1 <= numero4(contador);
		elsif destruidos/100 = 5 then
			color_numero1 <= numero5(contador);
		elsif destruidos/100 = 6 then
			color_numero1 <= numero6(contador);
		elsif destruidos/100 = 7 then
			color_numero1 <= numero7(contador);
		elsif destruidos/100 = 8 then
			color_numero1 <= numero8(contador);
		elsif destruidos/100 = 9 then
			color_numero1 <= numero9(contador);
		end if;
	end process contador_numero1;
	--
	
	contador_numero2 : process (clk_vga, num2_vali) is
		variable contador : integer range -1 to 576 := -1;
	begin
		if rising_edge(clk_vga) then
			if num2_vali = '1' then
				contador := contador+1;
				if contador = 575 then
					contador := -1;
				end if;
			end if;
		end if;
		
		if (destruidos mod 100)/10 = 0 then
			color_numero2 <= numero0(contador);
		elsif (destruidos mod 100)/10 = 1 then
			color_numero2 <= numero1(contador);
		elsif (destruidos mod 100)/10 = 2 then
			color_numero2 <= numero2(contador);
		elsif (destruidos mod 100)/10 = 3 then
			color_numero2 <= numero3(contador);
		elsif (destruidos mod 100)/10 = 4 then
			color_numero2 <= numero4(contador);
		elsif (destruidos mod 100)/10 = 5 then
			color_numero2 <= numero5(contador);
		elsif (destruidos mod 100)/10 = 6 then
			color_numero2 <= numero6(contador);
		elsif (destruidos mod 100)/10 = 7 then
			color_numero2 <= numero7(contador);
		elsif (destruidos mod 100)/10 = 8 then
			color_numero2 <= numero8(contador);
		elsif (destruidos mod 100)/10 = 9 then
			color_numero2 <= numero9(contador);
		end if;
		
	end process contador_numero2;
	--
	
	contador_numero3 : process (clk_vga, num3_vali) is
		variable contador : integer range -1 to 576 := -1;
	begin
		if rising_edge(clk_vga) then
			if num3_vali = '1' then
				contador := contador+1;
				if contador = 575 then
					contador := -1;
				end if;
			end if;
		end if;
		
		if destruidos mod 10 = 0 then
			color_numero3 <= numero0(contador);
		elsif destruidos mod 10 = 1 then
			color_numero3 <= numero1(contador);
		elsif destruidos mod 10 = 2 then
			color_numero3 <= numero2(contador);
		elsif destruidos mod 10 = 3 then
			color_numero3 <= numero3(contador);
		elsif destruidos mod 10 = 4 then
			color_numero3 <= numero4(contador);
		elsif destruidos mod 10 = 5 then
			color_numero3 <= numero5(contador);
		elsif destruidos mod 10 = 6 then
			color_numero3 <= numero6(contador);
		elsif destruidos mod 10 = 7 then
			color_numero3 <= numero7(contador);
		elsif destruidos mod 10 = 8 then
			color_numero3 <= numero8(contador);
		elsif destruidos mod 10 = 9 then
			color_numero3 <= numero9(contador);
		end if;
	
	end process contador_numero3;
	--
	
	contador_cora1 : process (clk_vga, cor1_vali) is
		variable contador : integer range -1 to 576 := -1;
	begin
		if rising_edge(clk_vga) then
			if cor1_vali = '1' then
				contador := contador+1;
				if contador = 575 then
					contador := -1;
				end if;
			end if;
		end if;
		color_cora1 <= cora(contador);
	end process contador_cora1;
	--
	
	contador_cora2 : process (clk_vga, cor2_vali) is
		variable contador : integer range -1 to 576 := -1;
	begin
		if rising_edge(clk_vga) then
			if cor2_vali = '1' then
				contador := contador+1;
				if contador = 575 then
					contador := -1;
				end if;
			end if;
		end if;
		color_cora2 <= cora(contador);
	end process contador_cora2;
	--
	
	contador_cora3 : process (clk_vga, cor3_vali) is
		variable contador : integer range -1 to 576 := -1;
	begin
		if rising_edge(clk_vga) then
			if cor3_vali = '1' then
				contador := contador+1;
				if contador = 575 then
					contador := -1;
				end if;
			end if;
		end if;
		color_cora3 <= cora(contador);
	end process contador_cora3;
	--
	
	-- Proceso para mostrar en la pantalla el pixel que queremos con el color deseado
	mostrar_pixel:	process (clk_vga,pintar,color_nave,asteroide_valido) is
	begin
		if rising_edge(clk_vga) then
			if pintar = '1' then
				
				if nave_vali = '1' and color_nave /= x"000" then
						vga_color <= color_nave;
					
				elsif asteroide_valido = '1' then
					vga_color <= x"C82";
					
				elsif disparo_vali = '1' then
					vga_color <= x"F00";
				
				elsif num1_vali = '1' then
					vga_color <= color_numero1;
				
				elsif num2_vali = '1' then
					vga_color <= color_numero2;
				
				elsif num3_vali = '1' then
					vga_color <= color_numero3;
				
				elsif cor1_vali = '1' then
					vga_color <= color_cora1;
					
				elsif cor2_vali = '1' then
					vga_color <= color_cora2;
					
				elsif cor3_vali = '1' then
					vga_color <= color_cora3;
					
				elsif over_vali = '1' then
					vga_color <= color_over;
					
				else
					vga_color <= x"000";
				end if;
			end if;	
		end if;
	end process mostrar_pixel;
	--
	
	--nave_vali <= '1' when (column > despX and column < despX+tam+1 and row > despY and row < despY+tam+1) else '0';
	nave_vali <= '1' when (column > despX and column < despX+tam+1 and row > v_video-tam-1 and row <= v_video-1) else '0';
	over_vali <= '1' when (vidas = 0 and column > 270 and column < 371 and row > 190 and row < 291) else '0';
	
	-- Definimos los asteroides que apareceran en la pantalla
	ast_vali0 <= '1' when ((row-desp_asteroide0)**2 + (column-posX_asteroide0)**2 < radio_asteroide**2) else '0';
	ast_vali1 <= '1' when ((row-desp_asteroide1)**2 + (column-posX_asteroide1)**2 < radio_asteroide**2) else '0';
	ast_vali2 <= '1' when ((row-desp_asteroide2)**2 + (column-posX_asteroide2)**2 < radio_asteroide**2) else '0';
	ast_vali3 <= '1' when ((row-desp_asteroide3)**2 + (column-posX_asteroide3)**2 < radio_asteroide**2) else '0';
	ast_vali4 <= '1' when ((row-desp_asteroide4)**2 + (column-posX_asteroide4)**2 < radio_asteroide**2) else '0';
	ast_vali5 <= '1' when ((row-desp_asteroide5)**2 + (column-posX_asteroide5)**2 < radio_asteroide**2) else '0';
	ast_vali6 <= '1' when ((row-desp_asteroide6)**2 + (column-posX_asteroide6)**2 < radio_asteroide**2) else '0';
	ast_vali7 <= '1' when ((row-desp_asteroide7)**2 + (column-posX_asteroide7)**2 < radio_asteroide**2) else '0';
	
	-- colorea disparo
	disparo_vali <= '1' when (recarga='0' and column > posx_disparo and column < posx_disparo+tam_disp+1 and row > desp_disparo and row < desp_disparo+tam_disp+1) else '0';
	
	--validaciones asteroide
	asteroide_valido <= ast_vali0 or ast_vali1 or ast_vali2 or ast_vali3 or ast_vali4 or ast_vali5 or ast_vali6 or ast_vali7;
	
	-- Validaciones para los numeros
	num1_vali <= '1' when (column>530 and column<555 and row>60 and row<85) else '0';
	num2_vali <= '1' when (column>555 and column<580 and row>60 and row<85) else '0';
	num3_vali <= '1' when (column>580 and column<605 and row>60 and row<85) else '0';
	
	-- Validaciones para mostrar los corazones de las vidas
	cor1_vali <= '1' when (vidas=3 and column>530 and column<555 and row>450 and row<475) else '0';
	cor2_vali <= '1' when (vidas>=2 and column>555 and column<580 and row>450 and row<475) else '0';
	cor3_vali <= '1' when (vidas>=1 and column>580 and column<605 and row>450 and row<475) else '0';
	
	vga_R <= vga_color(11 downto 8);
	vga_G <= vga_color(7 downto 4);
	vga_B <= vga_color(3 downto 0);
	
end architecture behavioral;